`include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype_FD.sv"

program automatic PATTERN(input clk, INF.PATTERN inf);
import usertype::*;

integer i;
Action now_action, previous_action;
Action action[400:0];
Restaurant_id res_id[400:0];
food_ID_servings food[400:0];
Delivery_man_id man_id[400:0];
Ctm_Info ctm[400:0];
Error_Msg message[400:0];
logic[63:0] answer[400:0];

initial begin
    inf.rst_n = 1;
    inf.act_valid = 0;
    inf.res_valid = 0;
    inf.food_valid = 0;
    inf.id_valid = 0;
    inf.cus_valid = 0;
    inf.D = 'bx;

    initial_action;
    initial_res;
    initial_food;
    initial_man;
    initial_ctm;
    initial_message;
    initial_answer;
    
    reset_task;

    previous_action = No_action;
    now_action = No_action;

    for(i = 1; i < 401; i = i + 1) begin 
        action_task;
        case(now_action)
            Take: begin 
                deliver_man_task;
                customer_task;
            end
            Deliver: begin
                deliver_man_task;
            end
            Order: begin 
                restaurant_task;
                food_task;
            end
            Cancel: begin 
                restaurant_task;
                food_task;
                deliver_man_task;
            end
        endcase
        wait_task;
        answer_task;
    end

    $finish;
end

task reset_task;
begin
    force clk = 0;
    #1 inf.rst_n = 0;
    #1 inf.rst_n = 1;
    #1 release clk;
end
endtask

task action_task;
begin 
    if(i === 87) begin 
        repeat(9) @(negedge clk);
    end
    else begin 
        repeat(1) @(negedge clk);
    end
    inf.act_valid = 1;
    previous_action = now_action;
    now_action = action[i];
    inf.D.d_act[0] = now_action;
    @(negedge clk);
    inf.act_valid = 0;
    inf.D = 'bx;
end
endtask

task restaurant_task;
begin 
    if(!(previous_action === Order && now_action === Order && res_id[i - 1] === res_id[i])) begin
        repeat(1) @(negedge clk);
        inf.res_valid = 1;
        inf.D.d_res_id[0] = res_id[i];
        @(negedge clk);
        inf.res_valid = 0;
        inf.D = 'bx;
    end
end
endtask

task food_task;
begin 
    if(i === 387) begin 
        repeat(5) @(negedge clk);
    end
    else begin 
        repeat(1) @(negedge clk);
    end
    inf.food_valid = 1;
    inf.D.d_food_ID_ser[0] = food[i];
    @(negedge clk);
    inf.food_valid = 0;
    inf.D = 'bx;
end
endtask

task deliver_man_task;
begin 
    if(!(previous_action === Take && now_action == Take && man_id[i - 1] === man_id[i])) begin
        repeat(1) @(negedge clk);
        inf.id_valid = 1;
        inf.D.d_id[0] = man_id[i];
        @(negedge clk);
        inf.id_valid = 0;
        inf.D = 'bx;
    end
end
endtask

task customer_task;
begin 
    repeat(1) @(negedge clk);
    inf.cus_valid = 1;
    inf.D.d_ctm_info[0] = ctm[i];
    @(negedge clk);
    inf.cus_valid = 0;
    inf.D = 'bx;
end
endtask

task wait_task;
begin 
    while(!inf.out_valid) @(negedge clk);
end
endtask

task answer_task;
begin 
    if(i > 200) begin 
        if(inf.out_info !== answer[i] || !inf.complete) begin 
            $display("Wrong Answer");
            $fatal;
        end
        else @(negedge clk);
    end
    else begin 
        if(inf.err_msg !== message[i] || inf.complete) begin 
            $display("Wrong Answer");
            $fatal;
        end
        else @(negedge clk);
    end
end
endtask

task initial_action;
begin
    action[  0] = No_action;
    action[  1] = Order;
    action[  2] = Take;
    action[  3] = Order;
    action[  4] = Take;
    action[  5] = Order;
    action[  6] = Take;
    action[  7] = Order;
    action[  8] = Take;
    action[  9] = Order;
    action[ 10] = Take;
    action[ 11] = Order;
    action[ 12] = Take;
    action[ 13] = Order;
    action[ 14] = Take;
    action[ 15] = Order;
    action[ 16] = Take;
    action[ 17] = Order;
    action[ 18] = Take;
    action[ 19] = Order;
    action[ 20] = Take;
    action[ 21] = Order;
    action[ 22] = Cancel;
    action[ 23] = Order;
    action[ 24] = Cancel;
    action[ 25] = Order;
    action[ 26] = Cancel;
    action[ 27] = Order;
    action[ 28] = Cancel;
    action[ 29] = Order;
    action[ 30] = Cancel;
    action[ 31] = Order;
    action[ 32] = Cancel;
    action[ 33] = Order;
    action[ 34] = Cancel;
    action[ 35] = Order;
    action[ 36] = Cancel;
    action[ 37] = Order;
    action[ 38] = Cancel;
    action[ 39] = Order;
    action[ 40] = Cancel;
    action[ 41] = Order;
    action[ 42] = Deliver;
    action[ 43] = Order;
    action[ 44] = Deliver;
    action[ 45] = Order;
    action[ 46] = Deliver;
    action[ 47] = Order;
    action[ 48] = Deliver;
    action[ 49] = Order;
    action[ 50] = Deliver;
    action[ 51] = Order;
    action[ 52] = Deliver;
    action[ 53] = Order;
    action[ 54] = Deliver;
    action[ 55] = Order;
    action[ 56] = Deliver;
    action[ 57] = Order;
    action[ 58] = Deliver;
    action[ 59] = Order;
    action[ 60] = Deliver;
    action[ 61] = Take;
    action[ 62] = Deliver;
    action[ 63] = Take;
    action[ 64] = Deliver;
    action[ 65] = Take;
    action[ 66] = Deliver;
    action[ 67] = Take;
    action[ 68] = Deliver;
    action[ 69] = Take;
    action[ 70] = Deliver;
    action[ 71] = Take;
    action[ 72] = Deliver;
    action[ 73] = Take;
    action[ 74] = Deliver;
    action[ 75] = Take;
    action[ 76] = Deliver;
    action[ 77] = Take;
    action[ 78] = Deliver;
    action[ 79] = Take;
    action[ 80] = Deliver;
    action[ 81] = Cancel;
    action[ 82] = Deliver;
    action[ 83] = Cancel;
    action[ 84] = Deliver;
    action[ 85] = Cancel;
    action[ 86] = Deliver;
    action[ 87] = Cancel;
    action[ 88] = Deliver;
    action[ 89] = Cancel;
    action[ 90] = Deliver;
    action[ 91] = Cancel;
    action[ 92] = Deliver;
    action[ 93] = Cancel;
    action[ 94] = Deliver;
    action[ 95] = Cancel;
    action[ 96] = Deliver;
    action[ 97] = Cancel;
    action[ 98] = Deliver;
    action[ 99] = Cancel;
    action[100] = Deliver;
    action[101] = Deliver;
    action[102] = Deliver;
    action[103] = Deliver;
    action[104] = Deliver;
    action[105] = Deliver;
    action[106] = Deliver;
    action[107] = Deliver;
    action[108] = Deliver;
    action[109] = Deliver;
    action[110] = Deliver;
    action[111] = Cancel;
    action[112] = Cancel;
    action[113] = Cancel;
    action[114] = Cancel;
    action[115] = Cancel;
    action[116] = Cancel;
    action[117] = Cancel;
    action[118] = Cancel;
    action[119] = Cancel;
    action[120] = Cancel;
    action[121] = Cancel;
    action[122] = Cancel;
    action[123] = Cancel;
    action[124] = Cancel;
    action[125] = Cancel;
    action[126] = Cancel;
    action[127] = Cancel;
    action[128] = Cancel;
    action[129] = Cancel;
    action[130] = Cancel;
    action[131] = Cancel;
    action[132] = Cancel;
    action[133] = Cancel;
    action[134] = Cancel;
    action[135] = Cancel;
    action[136] = Cancel;
    action[137] = Cancel;
    action[138] = Cancel;
    action[139] = Cancel;
    action[140] = Cancel;
    action[141] = Cancel;
    action[142] = Cancel;
    action[143] = Cancel;
    action[144] = Cancel;
    action[145] = Cancel;
    action[146] = Cancel;
    action[147] = Cancel;
    action[148] = Cancel;
    action[149] = Cancel;
    action[150] = Cancel;
    action[151] = Take;
    action[152] = Cancel;
    action[153] = Take;
    action[154] = Cancel;
    action[155] = Take;
    action[156] = Cancel;
    action[157] = Take;
    action[158] = Cancel;
    action[159] = Take;
    action[160] = Cancel;
    action[161] = Take;
    action[162] = Cancel;
    action[163] = Take;
    action[164] = Cancel;
    action[165] = Take;
    action[166] = Cancel;
    action[167] = Take;
    action[168] = Cancel;
    action[169] = Take;
    action[170] = Cancel;
    action[171] = Take;
    action[172] = Take;
    action[173] = Take;
    action[174] = Take;
    action[175] = Take;
    action[176] = Take;
    action[177] = Take;
    action[178] = Take;
    action[179] = Take;
    action[180] = Take;
    action[181] = Take;
    action[182] = Take;
    action[183] = Take;
    action[184] = Take;
    action[185] = Take;
    action[186] = Take;
    action[187] = Take;
    action[188] = Take;
    action[189] = Take;
    action[190] = Take;
    action[191] = Take;
    action[192] = Take;
    action[193] = Take;
    action[194] = Take;
    action[195] = Take;
    action[196] = Take;
    action[197] = Take;
    action[198] = Take;
    action[199] = Take;
    action[200] = Take;
    action[201] = Deliver;
    action[202] = Deliver;
    action[203] = Deliver;
    action[204] = Deliver;
    action[205] = Deliver;
    action[206] = Deliver;
    action[207] = Deliver;
    action[208] = Deliver;
    action[209] = Deliver;
    action[210] = Deliver;
    action[211] = Deliver;
    action[212] = Deliver;
    action[213] = Deliver;
    action[214] = Deliver;
    action[215] = Deliver;
    action[216] = Deliver;
    action[217] = Deliver;
    action[218] = Deliver;
    action[219] = Deliver;
    action[220] = Deliver;
    action[221] = Deliver;
    action[222] = Deliver;
    action[223] = Deliver;
    action[224] = Deliver;
    action[225] = Deliver;
    action[226] = Deliver;
    action[227] = Deliver;
    action[228] = Deliver;
    action[229] = Deliver;
    action[230] = Deliver;
    action[231] = Deliver;
    action[232] = Deliver;
    action[233] = Deliver;
    action[234] = Deliver;
    action[235] = Deliver;
    action[236] = Deliver;
    action[237] = Deliver;
    action[238] = Deliver;
    action[239] = Deliver;
    action[240] = Deliver;
    action[241] = Deliver;
    action[242] = Deliver;
    action[243] = Deliver;
    action[244] = Deliver;
    action[245] = Deliver;
    action[246] = Deliver;
    action[247] = Deliver;
    action[248] = Deliver;
    action[249] = Deliver;
    action[250] = Deliver;
    action[251] = Deliver;
    action[252] = Deliver;
    action[253] = Deliver;
    action[254] = Deliver;
    action[255] = Deliver;
    action[256] = Deliver;
    action[257] = Deliver;
    action[258] = Deliver;
    action[259] = Deliver;
    action[260] = Deliver;
    action[261] = Deliver;
    action[262] = Deliver;
    action[263] = Deliver;
    action[264] = Deliver;
    action[265] = Deliver;
    action[266] = Deliver;
    action[267] = Deliver;
    action[268] = Deliver;
    action[269] = Deliver;
    action[270] = Deliver;
    action[271] = Deliver;
    action[272] = Deliver;
    action[273] = Deliver;
    action[274] = Deliver;
    action[275] = Deliver;
    action[276] = Deliver;
    action[277] = Deliver;
    action[278] = Deliver;
    action[279] = Deliver;
    action[280] = Deliver;
    action[281] = Deliver;
    action[282] = Deliver;
    action[283] = Deliver;
    action[284] = Deliver;
    action[285] = Deliver;
    action[286] = Deliver;
    action[287] = Order;
    action[288] = Order;
    action[289] = Order;
    action[290] = Order;
    action[291] = Order;
    action[292] = Order;
    action[293] = Order;
    action[294] = Order;
    action[295] = Order;
    action[296] = Order;
    action[297] = Order;
    action[298] = Order;
    action[299] = Order;
    action[300] = Order;
    action[301] = Order;
    action[302] = Order;
    action[303] = Order;
    action[304] = Order;
    action[305] = Order;
    action[306] = Order;
    action[307] = Order;
    action[308] = Order;
    action[309] = Order;
    action[310] = Order;
    action[311] = Order;
    action[312] = Order;
    action[313] = Order;
    action[314] = Order;
    action[315] = Order;
    action[316] = Order;
    action[317] = Order;
    action[318] = Order;
    action[319] = Order;
    action[320] = Order;
    action[321] = Order;
    action[322] = Order;
    action[323] = Order;
    action[324] = Order;
    action[325] = Order;
    action[326] = Order;
    action[327] = Order;
    action[328] = Order;
    action[329] = Order;
    action[330] = Order;
    action[331] = Order;
    action[332] = Order;
    action[333] = Order;
    action[334] = Order;
    action[335] = Order;
    action[336] = Order;
    action[337] = Order;
    action[338] = Order;
    action[339] = Order;
    action[340] = Order;
    action[341] = Order;
    action[342] = Order;
    action[343] = Order;
    action[344] = Order;
    action[345] = Order;
    action[346] = Order;
    action[347] = Order;
    action[348] = Order;
    action[349] = Order;
    action[350] = Order;
    action[351] = Order;
    action[352] = Order;
    action[353] = Order;
    action[354] = Order;
    action[355] = Order;
    action[356] = Order;
    action[357] = Order;
    action[358] = Order;
    action[359] = Order;
    action[360] = Order;
    action[361] = Order;
    action[362] = Order;
    action[363] = Order;
    action[364] = Order;
    action[365] = Order;
    action[366] = Order;
    action[367] = Order;
    action[368] = Order;
    action[369] = Order;
    action[370] = Order;
    action[371] = Order;
    action[372] = Order;
    action[373] = Order;
    action[374] = Order;
    action[375] = Order;
    action[376] = Order;
    action[377] = Order;
    action[378] = Order;
    action[379] = Order;
    action[380] = Order;
    action[381] = Order;
    action[382] = Order;
    action[383] = Order;
    action[384] = Order;
    action[385] = Order;
    action[386] = Order;
    action[387] = Order;
    action[388] = Order;
    action[389] = Order;
    action[390] = Order;
    action[391] = Order;
    action[392] = Order;
    action[393] = Order;
    action[394] = Order;
    action[395] = Cancel;
    action[396] = Take;
    action[397] = Take;
    action[398] = Cancel;
    action[399] = Cancel;
    action[400] = Cancel;
end
endtask

task initial_res;
begin
    res_id[  0] = 0;
    res_id[  1] = 254;
    res_id[  2] = 0;
    res_id[  3] = 0;
    res_id[  4] = 0;
    res_id[  5] = 0;
    res_id[  6] = 0;
    res_id[  7] = 0;
    res_id[  8] = 0;
    res_id[  9] = 0;
    res_id[ 10] = 0;
    res_id[ 11] = 0;
    res_id[ 12] = 0;
    res_id[ 13] = 0;
    res_id[ 14] = 0;
    res_id[ 15] = 0;
    res_id[ 16] = 0;
    res_id[ 17] = 0;
    res_id[ 18] = 0;
    res_id[ 19] = 0;
    res_id[ 20] = 0;
    res_id[ 21] = 0;
    res_id[ 22] = 0;
    res_id[ 23] = 0;
    res_id[ 24] = 0;
    res_id[ 25] = 0;
    res_id[ 26] = 0;
    res_id[ 27] = 0;
    res_id[ 28] = 0;
    res_id[ 29] = 0;
    res_id[ 30] = 0;
    res_id[ 31] = 0;
    res_id[ 32] = 0;
    res_id[ 33] = 0;
    res_id[ 34] = 0;
    res_id[ 35] = 0;
    res_id[ 36] = 0;
    res_id[ 37] = 0;
    res_id[ 38] = 0;
    res_id[ 39] = 0;
    res_id[ 40] = 0;
    res_id[ 41] = 0;
    res_id[ 42] = 0;
    res_id[ 43] = 0;
    res_id[ 44] = 0;
    res_id[ 45] = 0;
    res_id[ 46] = 0;
    res_id[ 47] = 0;
    res_id[ 48] = 0;
    res_id[ 49] = 0;
    res_id[ 50] = 0;
    res_id[ 51] = 0;
    res_id[ 52] = 0;
    res_id[ 53] = 0;
    res_id[ 54] = 0;
    res_id[ 55] = 0;
    res_id[ 56] = 0;
    res_id[ 57] = 0;
    res_id[ 58] = 0;
    res_id[ 59] = 0;
    res_id[ 60] = 0;
    res_id[ 61] = 0;
    res_id[ 62] = 0;
    res_id[ 63] = 0;
    res_id[ 64] = 0;
    res_id[ 65] = 0;
    res_id[ 66] = 0;
    res_id[ 67] = 0;
    res_id[ 68] = 0;
    res_id[ 69] = 0;
    res_id[ 70] = 0;
    res_id[ 71] = 0;
    res_id[ 72] = 0;
    res_id[ 73] = 0;
    res_id[ 74] = 0;
    res_id[ 75] = 0;
    res_id[ 76] = 0;
    res_id[ 77] = 0;
    res_id[ 78] = 0;
    res_id[ 79] = 0;
    res_id[ 80] = 0;
    res_id[ 81] = 0;
    res_id[ 82] = 0;
    res_id[ 83] = 0;
    res_id[ 84] = 0;
    res_id[ 85] = 0;
    res_id[ 86] = 0;
    res_id[ 87] = 0;
    res_id[ 88] = 0;
    res_id[ 89] = 0;
    res_id[ 90] = 0;
    res_id[ 91] = 0;
    res_id[ 92] = 0;
    res_id[ 93] = 0;
    res_id[ 94] = 0;
    res_id[ 95] = 0;
    res_id[ 96] = 0;
    res_id[ 97] = 0;
    res_id[ 98] = 0;
    res_id[ 99] = 0;
    res_id[100] = 0;
    res_id[101] = 0;
    res_id[102] = 0;
    res_id[103] = 0;
    res_id[104] = 0;
    res_id[105] = 0;
    res_id[106] = 0;
    res_id[107] = 0;
    res_id[108] = 0;
    res_id[109] = 0;
    res_id[110] = 0;
    res_id[111] = 0;
    res_id[112] = 0;
    res_id[113] = 0;
    res_id[114] = 0;
    res_id[115] = 0;
    res_id[116] = 0;
    res_id[117] = 0;
    res_id[118] = 0;
    res_id[119] = 0;
    res_id[120] = 0;
    res_id[121] = 0;
    res_id[122] = 0;
    res_id[123] = 0;
    res_id[124] = 0;
    res_id[125] = 0;
    res_id[126] = 0;
    res_id[127] = 0;
    res_id[128] = 0;
    res_id[129] = 0;
    res_id[130] = 0;
    res_id[131] = 0;
    res_id[132] = 0;
    res_id[133] = 0;
    res_id[134] = 0;
    res_id[135] = 0;
    res_id[136] = 0;
    res_id[137] = 0;
    res_id[138] = 0;
    res_id[139] = 0;
    res_id[140] = 0;
    res_id[141] = 255;
    res_id[142] = 255;
    res_id[143] = 0;
    res_id[144] = 255;
    res_id[145] = 0;
    res_id[146] = 255;
    res_id[147] = 255;
    res_id[148] = 255;
    res_id[149] = 255;
    res_id[150] = 255;
    res_id[151] = 0;
    res_id[152] = 255;
    res_id[153] = 0;
    res_id[154] = 255;
    res_id[155] = 0;
    res_id[156] = 255;
    res_id[157] = 0;
    res_id[158] = 255;
    res_id[159] = 0;
    res_id[160] = 255;
    res_id[161] = 0;
    res_id[162] = 255;
    res_id[163] = 0;
    res_id[164] = 255;
    res_id[165] = 0;
    res_id[166] = 255;
    res_id[167] = 0;
    res_id[168] = 255;
    res_id[169] = 0;
    res_id[170] = 255;
    res_id[171] = 0;
    res_id[172] = 0;
    res_id[173] = 0;
    res_id[174] = 0;
    res_id[175] = 0;
    res_id[176] = 0;
    res_id[177] = 0;
    res_id[178] = 0;
    res_id[179] = 0;
    res_id[180] = 0;
    res_id[181] = 0;
    res_id[182] = 0;
    res_id[183] = 0;
    res_id[184] = 0;
    res_id[185] = 0;
    res_id[186] = 0;
    res_id[187] = 0;
    res_id[188] = 0;
    res_id[189] = 0;
    res_id[190] = 0;
    res_id[191] = 0;
    res_id[192] = 0;
    res_id[193] = 0;
    res_id[194] = 0;
    res_id[195] = 0;
    res_id[196] = 0;
    res_id[197] = 0;
    res_id[198] = 0;
    res_id[199] = 0;
    res_id[200] = 0;
    res_id[201] = 0;
    res_id[202] = 0;
    res_id[203] = 0;
    res_id[204] = 0;
    res_id[205] = 0;
    res_id[206] = 0;
    res_id[207] = 0;
    res_id[208] = 0;
    res_id[209] = 0;
    res_id[210] = 0;
    res_id[211] = 0;
    res_id[212] = 0;
    res_id[213] = 0;
    res_id[214] = 0;
    res_id[215] = 0;
    res_id[216] = 0;
    res_id[217] = 0;
    res_id[218] = 0;
    res_id[219] = 0;
    res_id[220] = 0;
    res_id[221] = 0;
    res_id[222] = 0;
    res_id[223] = 0;
    res_id[224] = 0;
    res_id[225] = 0;
    res_id[226] = 0;
    res_id[227] = 0;
    res_id[228] = 0;
    res_id[229] = 0;
    res_id[230] = 0;
    res_id[231] = 0;
    res_id[232] = 0;
    res_id[233] = 0;
    res_id[234] = 0;
    res_id[235] = 0;
    res_id[236] = 0;
    res_id[237] = 0;
    res_id[238] = 0;
    res_id[239] = 0;
    res_id[240] = 0;
    res_id[241] = 0;
    res_id[242] = 0;
    res_id[243] = 0;
    res_id[244] = 0;
    res_id[245] = 0;
    res_id[246] = 0;
    res_id[247] = 0;
    res_id[248] = 0;
    res_id[249] = 0;
    res_id[250] = 0;
    res_id[251] = 0;
    res_id[252] = 0;
    res_id[253] = 0;
    res_id[254] = 0;
    res_id[255] = 0;
    res_id[256] = 0;
    res_id[257] = 0;
    res_id[258] = 0;
    res_id[259] = 0;
    res_id[260] = 0;
    res_id[261] = 0;
    res_id[262] = 0;
    res_id[263] = 0;
    res_id[264] = 0;
    res_id[265] = 0;
    res_id[266] = 0;
    res_id[267] = 0;
    res_id[268] = 0;
    res_id[269] = 0;
    res_id[270] = 0;
    res_id[271] = 0;
    res_id[272] = 0;
    res_id[273] = 0;
    res_id[274] = 0;
    res_id[275] = 0;
    res_id[276] = 0;
    res_id[277] = 0;
    res_id[278] = 0;
    res_id[279] = 0;
    res_id[280] = 0;
    res_id[281] = 0;
    res_id[282] = 0;
    res_id[283] = 0;
    res_id[284] = 0;
    res_id[285] = 0;
    res_id[286] = 0;
    res_id[287] = 255;
    res_id[288] = 255;
    res_id[289] = 255;
    res_id[290] = 255;
    res_id[291] = 255;
    res_id[292] = 255;
    res_id[293] = 255;
    res_id[294] = 255;
    res_id[295] = 255;
    res_id[296] = 255;
    res_id[297] = 255;
    res_id[298] = 255;
    res_id[299] = 255;
    res_id[300] = 255;
    res_id[301] = 255;
    res_id[302] = 255;
    res_id[303] = 255;
    res_id[304] = 255;
    res_id[305] = 255;
    res_id[306] = 255;
    res_id[307] = 255;
    res_id[308] = 255;
    res_id[309] = 255;
    res_id[310] = 255;
    res_id[311] = 255;
    res_id[312] = 255;
    res_id[313] = 255;
    res_id[314] = 255;
    res_id[315] = 255;
    res_id[316] = 255;
    res_id[317] = 255;
    res_id[318] = 255;
    res_id[319] = 255;
    res_id[320] = 255;
    res_id[321] = 255;
    res_id[322] = 255;
    res_id[323] = 255;
    res_id[324] = 255;
    res_id[325] = 255;
    res_id[326] = 255;
    res_id[327] = 255;
    res_id[328] = 255;
    res_id[329] = 255;
    res_id[330] = 255;
    res_id[331] = 255;
    res_id[332] = 255;
    res_id[333] = 255;
    res_id[334] = 255;
    res_id[335] = 255;
    res_id[336] = 255;
    res_id[337] = 255;
    res_id[338] = 255;
    res_id[339] = 255;
    res_id[340] = 255;
    res_id[341] = 255;
    res_id[342] = 255;
    res_id[343] = 255;
    res_id[344] = 255;
    res_id[345] = 255;
    res_id[346] = 255;
    res_id[347] = 255;
    res_id[348] = 255;
    res_id[349] = 255;
    res_id[350] = 255;
    res_id[351] = 255;
    res_id[352] = 255;
    res_id[353] = 255;
    res_id[354] = 255;
    res_id[355] = 255;
    res_id[356] = 255;
    res_id[357] = 255;
    res_id[358] = 255;
    res_id[359] = 255;
    res_id[360] = 255;
    res_id[361] = 255;
    res_id[362] = 255;
    res_id[363] = 255;
    res_id[364] = 255;
    res_id[365] = 255;
    res_id[366] = 255;
    res_id[367] = 255;
    res_id[368] = 255;
    res_id[369] = 255;
    res_id[370] = 255;
    res_id[371] = 255;
    res_id[372] = 255;
    res_id[373] = 255;
    res_id[374] = 255;
    res_id[375] = 255;
    res_id[376] = 255;
    res_id[377] = 255;
    res_id[378] = 255;
    res_id[379] = 255;
    res_id[380] = 255;
    res_id[381] = 255;
    res_id[382] = 255;
    res_id[383] = 255;
    res_id[384] = 255;
    res_id[385] = 255;
    res_id[386] = 255;
    res_id[387] = 255;
    res_id[388] = 255;
    res_id[389] = 255;
    res_id[390] = 255;
    res_id[391] = 255;
    res_id[392] = 255;
    res_id[393] = 255;
    res_id[394] = 255;
    res_id[395] = 255;
    res_id[396] = 255;
    res_id[397] = 255;
    res_id[398] = 1;
    res_id[399] = 255;
    res_id[400] = 255;
end
endtask

task initial_food;
begin
    food[  0] = 6'b0;
    food[  1] = 6'h3f;
    food[  2] = 6'b0;
    food[  3] = 6'h3f;
    food[  4] = 6'b0;
    food[  5] = 6'h3f;
    food[  6] = 6'b0;
    food[  7] = 6'h3f;
    food[  8] = 6'b0;
    food[  9] = 6'h3f;
    food[ 10] = 6'b0;
    food[ 11] = 6'h3f;
    food[ 12] = 6'b0;
    food[ 13] = 6'h3f;
    food[ 14] = 6'b0;
    food[ 15] = 6'h3f;
    food[ 16] = 6'b0;
    food[ 17] = 6'h3f;
    food[ 18] = 6'b0;
    food[ 19] = 6'h3f;
    food[ 20] = 6'b0;
    food[ 21] = 6'h3f;
    food[ 22] = 6'h30;
    food[ 23] = 6'h3f;
    food[ 24] = 6'h30;
    food[ 25] = 6'h3f;
    food[ 26] = 6'h30;
    food[ 27] = 6'h3f;
    food[ 28] = 6'h30;
    food[ 29] = 6'h3f;
    food[ 30] = 6'h30;
    food[ 31] = 6'h3f;
    food[ 32] = 6'h30;
    food[ 33] = 6'h3f;
    food[ 34] = 6'h30;
    food[ 35] = 6'h3f;
    food[ 36] = 6'h30;
    food[ 37] = 6'h3f;
    food[ 38] = 6'h30;
    food[ 39] = 6'h3f;
    food[ 40] = 6'h30;
    food[ 41] = 6'h3f;
    food[ 42] = 6'b0;
    food[ 43] = 6'h3f;
    food[ 44] = 6'b0;
    food[ 45] = 6'h3f;
    food[ 46] = 6'b0;
    food[ 47] = 6'h3f;
    food[ 48] = 6'b0;
    food[ 49] = 6'h3f;
    food[ 50] = 6'b0;
    food[ 51] = 6'h3f;
    food[ 52] = 6'b0;
    food[ 53] = 6'h3f;
    food[ 54] = 6'b0;
    food[ 55] = 6'h3f;
    food[ 56] = 6'b0;
    food[ 57] = 6'h3f;
    food[ 58] = 6'b0;
    food[ 59] = 6'h3f;
    food[ 60] = 6'b0;
    food[ 61] = 6'b0;
    food[ 62] = 6'b0;
    food[ 63] = 6'b0;
    food[ 64] = 6'b0;
    food[ 65] = 6'b0;
    food[ 66] = 6'b0;
    food[ 67] = 6'b0;
    food[ 68] = 6'b0;
    food[ 69] = 6'b0;
    food[ 70] = 6'b0;
    food[ 71] = 6'b0;
    food[ 72] = 6'b0;
    food[ 73] = 6'b0;
    food[ 74] = 6'b0;
    food[ 75] = 6'b0;
    food[ 76] = 6'b0;
    food[ 77] = 6'b0;
    food[ 78] = 6'b0;
    food[ 79] = 6'b0;
    food[ 80] = 6'b0;
    food[ 81] = 6'h30;
    food[ 82] = 6'b0;
    food[ 83] = 6'h30;
    food[ 84] = 6'b0;
    food[ 85] = 6'h30;
    food[ 86] = 6'b0;
    food[ 87] = 6'h30;
    food[ 88] = 6'b0;
    food[ 89] = 6'h30;
    food[ 90] = 6'b0;
    food[ 91] = 6'h30;
    food[ 92] = 6'b0;
    food[ 93] = 6'h30;
    food[ 94] = 6'b0;
    food[ 95] = 6'h30;
    food[ 96] = 6'b0;
    food[ 97] = 6'h30;
    food[ 98] = 6'b0;
    food[ 99] = 6'h30;
    food[100] = 6'b0;
    food[101] = 6'b0;
    food[102] = 6'b0;
    food[103] = 6'b0;
    food[104] = 6'b0;
    food[105] = 6'b0;
    food[106] = 6'b0;
    food[107] = 6'b0;
    food[108] = 6'b0;
    food[109] = 6'b0;
    food[110] = 6'b0;
    food[111] = 6'h30;
    food[112] = 6'h30;
    food[113] = 6'h30;
    food[114] = 6'h30;
    food[115] = 6'h30;
    food[116] = 6'h30;
    food[117] = 6'h30;
    food[118] = 6'h30;
    food[119] = 6'h30;
    food[120] = 6'h30;
    food[121] = 6'h30;
    food[122] = 6'h30;
    food[123] = 6'h30;
    food[124] = 6'h30;
    food[125] = 6'h30;
    food[126] = 6'h30;
    food[127] = 6'h30;
    food[128] = 6'h30;
    food[129] = 6'h30;
    food[130] = 6'h30;
    food[131] = 6'h30;
    food[132] = 6'h30;
    food[133] = 6'h30;
    food[134] = 6'h30;
    food[135] = 6'h30;
    food[136] = 6'h30;
    food[137] = 6'h30;
    food[138] = 6'h30;
    food[139] = 6'h30;
    food[140] = 6'h30;
    food[141] = 6'h10;
    food[142] = 6'h10;
    food[143] = 6'h10;
    food[144] = 6'h10;
    food[145] = 6'h10;
    food[146] = 6'h10;
    food[147] = 6'h10;
    food[148] = 6'h10;
    food[149] = 6'h10;
    food[150] = 6'h10;
    food[151] = 6'b0;
    food[152] = 6'h10;
    food[153] = 6'b0;
    food[154] = 6'h10;
    food[155] = 6'b0;
    food[156] = 6'h10;
    food[157] = 6'b0;
    food[158] = 6'h10;
    food[159] = 6'b0;
    food[160] = 6'h10;
    food[161] = 6'b0;
    food[162] = 6'h10;
    food[163] = 6'b0;
    food[164] = 6'h10;
    food[165] = 6'b0;
    food[166] = 6'h10;
    food[167] = 6'b0;
    food[168] = 6'h10;
    food[169] = 6'b0;
    food[170] = 6'h10;
    food[171] = 6'b0;
    food[172] = 6'b0;
    food[173] = 6'b0;
    food[174] = 6'b0;
    food[175] = 6'b0;
    food[176] = 6'b0;
    food[177] = 6'b0;
    food[178] = 6'b0;
    food[179] = 6'b0;
    food[180] = 6'b0;
    food[181] = 6'b0;
    food[182] = 6'b0;
    food[183] = 6'b0;
    food[184] = 6'b0;
    food[185] = 6'b0;
    food[186] = 6'b0;
    food[187] = 6'b0;
    food[188] = 6'b0;
    food[189] = 6'b0;
    food[190] = 6'b0;
    food[191] = 6'b0;
    food[192] = 6'b0;
    food[193] = 6'b0;
    food[194] = 6'b0;
    food[195] = 6'b0;
    food[196] = 6'b0;
    food[197] = 6'b0;
    food[198] = 6'b0;
    food[199] = 6'b0;
    food[200] = 6'b0;
    food[201] = 6'b0;
    food[202] = 6'b0;
    food[203] = 6'b0;
    food[204] = 6'b0;
    food[205] = 6'b0;
    food[206] = 6'b0;
    food[207] = 6'b0;
    food[208] = 6'b0;
    food[209] = 6'b0;
    food[210] = 6'b0;
    food[211] = 6'b0;
    food[212] = 6'b0;
    food[213] = 6'b0;
    food[214] = 6'b0;
    food[215] = 6'b0;
    food[216] = 6'b0;
    food[217] = 6'b0;
    food[218] = 6'b0;
    food[219] = 6'b0;
    food[220] = 6'b0;
    food[221] = 6'b0;
    food[222] = 6'b0;
    food[223] = 6'b0;
    food[224] = 6'b0;
    food[225] = 6'b0;
    food[226] = 6'b0;
    food[227] = 6'b0;
    food[228] = 6'b0;
    food[229] = 6'b0;
    food[230] = 6'b0;
    food[231] = 6'b0;
    food[232] = 6'b0;
    food[233] = 6'b0;
    food[234] = 6'b0;
    food[235] = 6'b0;
    food[236] = 6'b0;
    food[237] = 6'b0;
    food[238] = 6'b0;
    food[239] = 6'b0;
    food[240] = 6'b0;
    food[241] = 6'b0;
    food[242] = 6'b0;
    food[243] = 6'b0;
    food[244] = 6'b0;
    food[245] = 6'b0;
    food[246] = 6'b0;
    food[247] = 6'b0;
    food[248] = 6'b0;
    food[249] = 6'b0;
    food[250] = 6'b0;
    food[251] = 6'b0;
    food[252] = 6'b0;
    food[253] = 6'b0;
    food[254] = 6'b0;
    food[255] = 6'b0;
    food[256] = 6'b0;
    food[257] = 6'b0;
    food[258] = 6'b0;
    food[259] = 6'b0;
    food[260] = 6'b0;
    food[261] = 6'b0;
    food[262] = 6'b0;
    food[263] = 6'b0;
    food[264] = 6'b0;
    food[265] = 6'b0;
    food[266] = 6'b0;
    food[267] = 6'b0;
    food[268] = 6'b0;
    food[269] = 6'b0;
    food[270] = 6'b0;
    food[271] = 6'b0;
    food[272] = 6'b0;
    food[273] = 6'b0;
    food[274] = 6'b0;
    food[275] = 6'b0;
    food[276] = 6'b0;
    food[277] = 6'b0;
    food[278] = 6'b0;
    food[279] = 6'b0;
    food[280] = 6'b0;
    food[281] = 6'b0;
    food[282] = 6'b0;
    food[283] = 6'b0;
    food[284] = 6'b0;
    food[285] = 6'b0;
    food[286] = 6'b0;
    food[287] = 6'h11;
    food[288] = 6'h11;
    food[289] = 6'h11;
    food[290] = 6'h11;
    food[291] = 6'h11;
    food[292] = 6'h11;
    food[293] = 6'h11;
    food[294] = 6'h11;
    food[295] = 6'h11;
    food[296] = 6'h11;
    food[297] = 6'h11;
    food[298] = 6'h11;
    food[299] = 6'h11;
    food[300] = 6'h11;
    food[301] = 6'h11;
    food[302] = 6'h11;
    food[303] = 6'h11;
    food[304] = 6'h11;
    food[305] = 6'h11;
    food[306] = 6'h11;
    food[307] = 6'h11;
    food[308] = 6'h11;
    food[309] = 6'h11;
    food[310] = 6'h11;
    food[311] = 6'h11;
    food[312] = 6'h11;
    food[313] = 6'h11;
    food[314] = 6'h11;
    food[315] = 6'h11;
    food[316] = 6'h11;
    food[317] = 6'h11;
    food[318] = 6'h11;
    food[319] = 6'h11;
    food[320] = 6'h11;
    food[321] = 6'h11;
    food[322] = 6'h11;
    food[323] = 6'h11;
    food[324] = 6'h11;
    food[325] = 6'h11;
    food[326] = 6'h11;
    food[327] = 6'h11;
    food[328] = 6'h11;
    food[329] = 6'h11;
    food[330] = 6'h11;
    food[331] = 6'h11;
    food[332] = 6'h11;
    food[333] = 6'h11;
    food[334] = 6'h11;
    food[335] = 6'h11;
    food[336] = 6'h11;
    food[337] = 6'h11;
    food[338] = 6'h11;
    food[339] = 6'h11;
    food[340] = 6'h11;
    food[341] = 6'h11;
    food[342] = 6'h11;
    food[343] = 6'h11;
    food[344] = 6'h11;
    food[345] = 6'h11;
    food[346] = 6'h11;
    food[347] = 6'h11;
    food[348] = 6'h11;
    food[349] = 6'h11;
    food[350] = 6'h11;
    food[351] = 6'h11;
    food[352] = 6'h11;
    food[353] = 6'h11;
    food[354] = 6'h11;
    food[355] = 6'h11;
    food[356] = 6'h11;
    food[357] = 6'h11;
    food[358] = 6'h11;
    food[359] = 6'h11;
    food[360] = 6'h11;
    food[361] = 6'h11;
    food[362] = 6'h11;
    food[363] = 6'h11;
    food[364] = 6'h11;
    food[365] = 6'h11;
    food[366] = 6'h11;
    food[367] = 6'h11;
    food[368] = 6'h11;
    food[369] = 6'h11;
    food[370] = 6'h11;
    food[371] = 6'h11;
    food[372] = 6'h11;
    food[373] = 6'h11;
    food[374] = 6'h11;
    food[375] = 6'h11;
    food[376] = 6'h11;
    food[377] = 6'h11;
    food[378] = 6'h11;
    food[379] = 6'h11;
    food[380] = 6'h11;
    food[381] = 6'h11;
    food[382] = 6'h11;
    food[383] = 6'h11;
    food[384] = 6'h11;
    food[385] = 6'h11;
    food[386] = 6'h11;
    food[387] = 6'h11;
    food[388] = 6'h11;
    food[389] = 6'h11;
    food[390] = 6'h11;
    food[391] = 6'h11;
    food[392] = 6'h11;
    food[393] = 6'h11;
    food[394] = 6'h11;
    food[395] = 6'h30;
    food[396] = 6'h11;
    food[397] = 6'h11;
    food[398] = 6'h10;
    food[399] = 6'h30;
    food[400] = 6'h30;
end
endtask

task initial_man;
begin
    man_id[  0] = 0;
    man_id[  1] = 0;
    man_id[  2] = 0;
    man_id[  3] = 1;
    man_id[  4] = 1;
    man_id[  5] = 2;
    man_id[  6] = 2;
    man_id[  7] = 3;
    man_id[  8] = 3;
    man_id[  9] = 4;
    man_id[ 10] = 4;
    man_id[ 11] = 5;
    man_id[ 12] = 5;
    man_id[ 13] = 6;
    man_id[ 14] = 6;
    man_id[ 15] = 7;
    man_id[ 16] = 7;
    man_id[ 17] = 8;
    man_id[ 18] = 8;
    man_id[ 19] = 9;
    man_id[ 20] = 9;
    man_id[ 21] = 10;
    man_id[ 22] = 10;
    man_id[ 23] = 11;
    man_id[ 24] = 11;
    man_id[ 25] = 12;
    man_id[ 26] = 12;
    man_id[ 27] = 13;
    man_id[ 28] = 13;
    man_id[ 29] = 14;
    man_id[ 30] = 14;
    man_id[ 31] = 15;
    man_id[ 32] = 15;
    man_id[ 33] = 16;
    man_id[ 34] = 16;
    man_id[ 35] = 17;
    man_id[ 36] = 17;
    man_id[ 37] = 18;
    man_id[ 38] = 18;
    man_id[ 39] = 19;
    man_id[ 40] = 19;
    man_id[ 41] = 20;
    man_id[ 42] = 20;
    man_id[ 43] = 21;
    man_id[ 44] = 21;
    man_id[ 45] = 22;
    man_id[ 46] = 22;
    man_id[ 47] = 23;
    man_id[ 48] = 23;
    man_id[ 49] = 24;
    man_id[ 50] = 24;
    man_id[ 51] = 25;
    man_id[ 52] = 25;
    man_id[ 53] = 26;
    man_id[ 54] = 26;
    man_id[ 55] = 27;
    man_id[ 56] = 27;
    man_id[ 57] = 28;
    man_id[ 58] = 28;
    man_id[ 59] = 29;
    man_id[ 60] = 29;
    man_id[ 61] = 30;
    man_id[ 62] = 31;
    man_id[ 63] = 32;
    man_id[ 64] = 33;
    man_id[ 65] = 34;
    man_id[ 66] = 35;
    man_id[ 67] = 36;
    man_id[ 68] = 37;
    man_id[ 69] = 38;
    man_id[ 70] = 39;
    man_id[ 71] = 40;
    man_id[ 72] = 41;
    man_id[ 73] = 42;
    man_id[ 74] = 43;
    man_id[ 75] = 44;
    man_id[ 76] = 45;
    man_id[ 77] = 46;
    man_id[ 78] = 47;
    man_id[ 79] = 48;
    man_id[ 80] = 49;
    man_id[ 81] = 50;
    man_id[ 82] = 51;
    man_id[ 83] = 52;
    man_id[ 84] = 53;
    man_id[ 85] = 54;
    man_id[ 86] = 55;
    man_id[ 87] = 56;
    man_id[ 88] = 57;
    man_id[ 89] = 58;
    man_id[ 90] = 59;
    man_id[ 91] = 60;
    man_id[ 92] = 61;
    man_id[ 93] = 62;
    man_id[ 94] = 63;
    man_id[ 95] = 64;
    man_id[ 96] = 65;
    man_id[ 97] = 66;
    man_id[ 98] = 67;
    man_id[ 99] = 68;
    man_id[100] = 69;
    man_id[101] = 70;
    man_id[102] = 71;
    man_id[103] = 72;
    man_id[104] = 73;
    man_id[105] = 74;
    man_id[106] = 75;
    man_id[107] = 76;
    man_id[108] = 77;
    man_id[109] = 78;
    man_id[110] = 79;
    man_id[111] = 80;
    man_id[112] = 81;
    man_id[113] = 82;
    man_id[114] = 83;
    man_id[115] = 84;
    man_id[116] = 85;
    man_id[117] = 86;
    man_id[118] = 87;
    man_id[119] = 88;
    man_id[120] = 89;
    man_id[121] = 90;
    man_id[122] = 91;
    man_id[123] = 92;
    man_id[124] = 93;
    man_id[125] = 94;
    man_id[126] = 95;
    man_id[127] = 96;
    man_id[128] = 97;
    man_id[129] = 98;
    man_id[130] = 99;
    man_id[131] = 100;
    man_id[132] = 101;
    man_id[133] = 102;
    man_id[134] = 103;
    man_id[135] = 104;
    man_id[136] = 105;
    man_id[137] = 106;
    man_id[138] = 107;
    man_id[139] = 108;
    man_id[140] = 109;
    man_id[141] = 110;
    man_id[142] = 111;
    man_id[143] = 112;
    man_id[144] = 113;
    man_id[145] = 114;
    man_id[146] = 115;
    man_id[147] = 116;
    man_id[148] = 117;
    man_id[149] = 118;
    man_id[150] = 119;
    man_id[151] = 120;
    man_id[152] = 121;
    man_id[153] = 122;
    man_id[154] = 123;
    man_id[155] = 124;
    man_id[156] = 125;
    man_id[157] = 126;
    man_id[158] = 127;
    man_id[159] = 128;
    man_id[160] = 129;
    man_id[161] = 130;
    man_id[162] = 131;
    man_id[163] = 132;
    man_id[164] = 133;
    man_id[165] = 134;
    man_id[166] = 135;
    man_id[167] = 136;
    man_id[168] = 137;
    man_id[169] = 138;
    man_id[170] = 139;
    man_id[171] = 140;
    man_id[172] = 141;
    man_id[173] = 142;
    man_id[174] = 143;
    man_id[175] = 144;
    man_id[176] = 145;
    man_id[177] = 146;
    man_id[178] = 147;
    man_id[179] = 148;
    man_id[180] = 149;
    man_id[181] = 150;
    man_id[182] = 151;
    man_id[183] = 152;
    man_id[184] = 153;
    man_id[185] = 154;
    man_id[186] = 155;
    man_id[187] = 156;
    man_id[188] = 157;
    man_id[189] = 158;
    man_id[190] = 159;
    man_id[191] = 160;
    man_id[192] = 161;
    man_id[193] = 162;
    man_id[194] = 163;
    man_id[195] = 164;
    man_id[196] = 165;
    man_id[197] = 166;
    man_id[198] = 167;
    man_id[199] = 168;
    man_id[200] = 169;
    man_id[201] = 170;
    man_id[202] = 171;
    man_id[203] = 172;
    man_id[204] = 173;
    man_id[205] = 174;
    man_id[206] = 175;
    man_id[207] = 176;
    man_id[208] = 177;
    man_id[209] = 178;
    man_id[210] = 179;
    man_id[211] = 180;
    man_id[212] = 181;
    man_id[213] = 182;
    man_id[214] = 183;
    man_id[215] = 184;
    man_id[216] = 185;
    man_id[217] = 186;
    man_id[218] = 187;
    man_id[219] = 188;
    man_id[220] = 189;
    man_id[221] = 190;
    man_id[222] = 191;
    man_id[223] = 192;
    man_id[224] = 193;
    man_id[225] = 194;
    man_id[226] = 195;
    man_id[227] = 196;
    man_id[228] = 197;
    man_id[229] = 198;
    man_id[230] = 199;
    man_id[231] = 200;
    man_id[232] = 201;
    man_id[233] = 202;
    man_id[234] = 203;
    man_id[235] = 204;
    man_id[236] = 205;
    man_id[237] = 206;
    man_id[238] = 207;
    man_id[239] = 208;
    man_id[240] = 209;
    man_id[241] = 210;
    man_id[242] = 211;
    man_id[243] = 212;
    man_id[244] = 213;
    man_id[245] = 214;
    man_id[246] = 215;
    man_id[247] = 216;
    man_id[248] = 217;
    man_id[249] = 218;
    man_id[250] = 219;
    man_id[251] = 220;
    man_id[252] = 221;
    man_id[253] = 222;
    man_id[254] = 223;
    man_id[255] = 224;
    man_id[256] = 225;
    man_id[257] = 226;
    man_id[258] = 227;
    man_id[259] = 228;
    man_id[260] = 229;
    man_id[261] = 230;
    man_id[262] = 231;
    man_id[263] = 232;
    man_id[264] = 233;
    man_id[265] = 234;
    man_id[266] = 235;
    man_id[267] = 236;
    man_id[268] = 237;
    man_id[269] = 238;
    man_id[270] = 239;
    man_id[271] = 240;
    man_id[272] = 241;
    man_id[273] = 242;
    man_id[274] = 243;
    man_id[275] = 244;
    man_id[276] = 245;
    man_id[277] = 246;
    man_id[278] = 247;
    man_id[279] = 248;
    man_id[280] = 249;
    man_id[281] = 250;
    man_id[282] = 251;
    man_id[283] = 252;
    man_id[284] = 253;
    man_id[285] = 254;
    man_id[286] = 255;
    man_id[287] = 0;
    man_id[288] = 0;
    man_id[289] = 0;
    man_id[290] = 0;
    man_id[291] = 0;
    man_id[292] = 0;
    man_id[293] = 0;
    man_id[294] = 0;
    man_id[295] = 0;
    man_id[296] = 0;
    man_id[297] = 0;
    man_id[298] = 0;
    man_id[299] = 0;
    man_id[300] = 0;
    man_id[301] = 0;
    man_id[302] = 0;
    man_id[303] = 0;
    man_id[304] = 0;
    man_id[305] = 0;
    man_id[306] = 0;
    man_id[307] = 0;
    man_id[308] = 0;
    man_id[309] = 0;
    man_id[310] = 0;
    man_id[311] = 0;
    man_id[312] = 0;
    man_id[313] = 0;
    man_id[314] = 0;
    man_id[315] = 0;
    man_id[316] = 0;
    man_id[317] = 0;
    man_id[318] = 0;
    man_id[319] = 0;
    man_id[320] = 0;
    man_id[321] = 0;
    man_id[322] = 0;
    man_id[323] = 0;
    man_id[324] = 0;
    man_id[325] = 0;
    man_id[326] = 0;
    man_id[327] = 0;
    man_id[328] = 0;
    man_id[329] = 0;
    man_id[330] = 0;
    man_id[331] = 0;
    man_id[332] = 0;
    man_id[333] = 0;
    man_id[334] = 0;
    man_id[335] = 0;
    man_id[336] = 0;
    man_id[337] = 0;
    man_id[338] = 0;
    man_id[339] = 0;
    man_id[340] = 0;
    man_id[341] = 0;
    man_id[342] = 0;
    man_id[343] = 0;
    man_id[344] = 0;
    man_id[345] = 0;
    man_id[346] = 0;
    man_id[347] = 0;
    man_id[348] = 0;
    man_id[349] = 0;
    man_id[350] = 0;
    man_id[351] = 0;
    man_id[352] = 0;
    man_id[353] = 0;
    man_id[354] = 0;
    man_id[355] = 0;
    man_id[356] = 0;
    man_id[357] = 0;
    man_id[358] = 0;
    man_id[359] = 0;
    man_id[360] = 0;
    man_id[361] = 0;
    man_id[362] = 0;
    man_id[363] = 0;
    man_id[364] = 0;
    man_id[365] = 0;
    man_id[366] = 0;
    man_id[367] = 0;
    man_id[368] = 0;
    man_id[369] = 0;
    man_id[370] = 0;
    man_id[371] = 0;
    man_id[372] = 0;
    man_id[373] = 0;
    man_id[374] = 0;
    man_id[375] = 0;
    man_id[376] = 0;
    man_id[377] = 0;
    man_id[378] = 0;
    man_id[379] = 0;
    man_id[380] = 0;
    man_id[381] = 0;
    man_id[382] = 0;
    man_id[383] = 0;
    man_id[384] = 0;
    man_id[385] = 0;
    man_id[386] = 0;
    man_id[387] = 0;
    man_id[388] = 0;
    man_id[389] = 0;
    man_id[390] = 0;
    man_id[391] = 0;
    man_id[392] = 0;
    man_id[393] = 0;
    man_id[394] = 0;
    man_id[395] = 168;
    man_id[396] = 1;
    man_id[397] = 1;
    man_id[398] = 1;
    man_id[399] = 169;
    man_id[400] = 170;
end
endtask

task initial_ctm;
begin
    ctm[ 20] = 16'h0000;
    ctm[  1] = 16'hffff;
    ctm[  2] = 16'hffff;
    ctm[  3] = 16'hffff;
    ctm[  4] = 16'hffff;
    ctm[  5] = 16'hffff;
    ctm[  6] = 16'hffff;
    ctm[  7] = 16'hffff;
    ctm[  8] = 16'hffff;
    ctm[  9] = 16'hffff;
    ctm[ 10] = 16'hffff;
    ctm[ 11] = 16'hffff;
    ctm[ 12] = 16'hffff;
    ctm[ 13] = 16'hffff;
    ctm[ 14] = 16'hffff;
    ctm[ 15] = 16'hffff;
    ctm[ 16] = 16'hffff;
    ctm[ 17] = 16'hffff;
    ctm[ 18] = 16'hffff;
    ctm[ 19] = 16'hffff;
    ctm[ 20] = 16'hffff;
    ctm[ 21] = 16'hffff;
    ctm[ 22] = 16'hffff;
    ctm[ 23] = 16'hffff;
    ctm[ 24] = 16'hffff;
    ctm[ 25] = 16'hffff;
    ctm[ 26] = 16'hffff;
    ctm[ 27] = 16'hffff;
    ctm[ 28] = 16'hffff;
    ctm[ 29] = 16'hffff;
    ctm[ 30] = 16'hffff;
    ctm[ 31] = 16'hffff;
    ctm[ 32] = 16'hffff;
    ctm[ 33] = 16'hffff;
    ctm[ 34] = 16'hffff;
    ctm[ 35] = 16'hffff;
    ctm[ 36] = 16'hffff;
    ctm[ 37] = 16'hffff;
    ctm[ 38] = 16'hffff;
    ctm[ 39] = 16'hffff;
    ctm[ 40] = 16'hffff;
    ctm[ 41] = 16'hffff;
    ctm[ 42] = 16'hffff;
    ctm[ 43] = 16'hffff;
    ctm[ 44] = 16'hffff;
    ctm[ 45] = 16'hffff;
    ctm[ 46] = 16'hffff;
    ctm[ 47] = 16'hffff;
    ctm[ 48] = 16'hffff;
    ctm[ 49] = 16'hffff;
    ctm[ 50] = 16'hffff;
    ctm[ 51] = 16'hffff;
    ctm[ 52] = 16'hffff;
    ctm[ 53] = 16'hffff;
    ctm[ 54] = 16'hffff;
    ctm[ 55] = 16'hffff;
    ctm[ 56] = 16'hffff;
    ctm[ 57] = 16'hffff;
    ctm[ 58] = 16'hffff;
    ctm[ 59] = 16'hffff;
    ctm[ 60] = 16'hffff;
    ctm[ 61] = 16'hffff;
    ctm[ 62] = 16'hffff;
    ctm[ 63] = 16'hffff;
    ctm[ 64] = 16'hffff;
    ctm[ 65] = 16'hffff;
    ctm[ 66] = 16'hffff;
    ctm[ 67] = 16'hffff;
    ctm[ 68] = 16'hffff;
    ctm[ 69] = 16'hffff;
    ctm[ 70] = 16'hffff;
    ctm[ 71] = 16'hffff;
    ctm[ 72] = 16'hffff;
    ctm[ 73] = 16'hffff;
    ctm[ 74] = 16'hffff;
    ctm[ 75] = 16'hffff;
    ctm[ 76] = 16'hffff;
    ctm[ 77] = 16'hffff;
    ctm[ 78] = 16'hffff;
    ctm[ 79] = 16'hffff;
    ctm[ 80] = 16'hffff;
    ctm[ 81] = 16'hffff;
    ctm[ 82] = 16'hffff;
    ctm[ 83] = 16'hffff;
    ctm[ 84] = 16'hffff;
    ctm[ 85] = 16'hffff;
    ctm[ 86] = 16'hffff;
    ctm[ 87] = 16'hffff;
    ctm[ 88] = 16'hffff;
    ctm[ 89] = 16'hffff;
    ctm[ 90] = 16'hffff;
    ctm[ 91] = 16'hffff;
    ctm[ 92] = 16'hffff;
    ctm[ 93] = 16'hffff;
    ctm[ 94] = 16'hffff;
    ctm[ 95] = 16'hffff;
    ctm[ 96] = 16'hffff;
    ctm[ 97] = 16'hffff;
    ctm[ 98] = 16'hffff;
    ctm[ 99] = 16'hffff;
    ctm[100] = 16'hffff;
    ctm[101] = 16'hffff;
    ctm[102] = 16'hffff;
    ctm[103] = 16'hffff;
    ctm[104] = 16'hffff;
    ctm[105] = 16'hffff;
    ctm[106] = 16'hffff;
    ctm[107] = 16'hffff;
    ctm[108] = 16'hffff;
    ctm[109] = 16'hffff;
    ctm[110] = 16'hffff;
    ctm[111] = 16'hffff;
    ctm[112] = 16'hffff;
    ctm[113] = 16'hffff;
    ctm[114] = 16'hffff;
    ctm[115] = 16'hffff;
    ctm[116] = 16'hffff;
    ctm[117] = 16'hffff;
    ctm[118] = 16'hffff;
    ctm[119] = 16'hffff;
    ctm[120] = 16'hffff;
    ctm[121] = 16'hffff;
    ctm[122] = 16'hffff;
    ctm[123] = 16'hffff;
    ctm[124] = 16'hffff;
    ctm[125] = 16'hffff;
    ctm[126] = 16'hffff;
    ctm[127] = 16'hffff;
    ctm[128] = 16'hffff;
    ctm[129] = 16'hffff;
    ctm[130] = 16'hffff;
    ctm[131] = 16'hffff;
    ctm[132] = 16'hffff;
    ctm[133] = 16'hffff;
    ctm[134] = 16'hffff;
    ctm[135] = 16'hffff;
    ctm[136] = 16'hffff;
    ctm[137] = 16'hffff;
    ctm[138] = 16'hffff;
    ctm[139] = 16'hffff;
    ctm[140] = 16'hffff;
    ctm[141] = 16'hffff;
    ctm[142] = 16'hffff;
    ctm[143] = 16'hffff;
    ctm[144] = 16'hffff;
    ctm[145] = 16'hffff;
    ctm[146] = 16'hffff;
    ctm[147] = 16'hffff;
    ctm[148] = 16'hffff;
    ctm[149] = 16'hffff;
    ctm[150] = 16'hffff;
    ctm[151] = 16'hffff;
    ctm[152] = 16'hffff;
    ctm[153] = 16'hffff;
    ctm[154] = 16'hffff;
    ctm[155] = 16'hffff;
    ctm[156] = 16'hffff;
    ctm[157] = 16'hffff;
    ctm[158] = 16'hffff;
    ctm[159] = 16'hffff;
    ctm[160] = 16'hffff;
    ctm[161] = 16'hffff;
    ctm[162] = 16'hffff;
    ctm[163] = 16'hffff;
    ctm[164] = 16'hffff;
    ctm[165] = 16'hffff;
    ctm[166] = 16'hffff;
    ctm[167] = 16'hffff;
    ctm[168] = 16'hffff;
    ctm[169] = 16'hffff;
    ctm[170] = 16'hffff;
    ctm[171] = 16'hffff;
    ctm[172] = 16'hffff;
    ctm[173] = 16'hffff;
    ctm[174] = 16'hffff;
    ctm[175] = 16'hffff;
    ctm[176] = 16'hffff;
    ctm[177] = 16'hffff;
    ctm[178] = 16'hffff;
    ctm[179] = 16'hffff;
    ctm[180] = 16'hffff;
    ctm[181] = 16'hffff;
    ctm[182] = 16'hffff;
    ctm[183] = 16'hffff;
    ctm[184] = 16'hffff;
    ctm[185] = 16'hffff;
    ctm[186] = 16'hffff;
    ctm[187] = 16'hffff;
    ctm[188] = 16'hffff;
    ctm[189] = 16'hffff;
    ctm[190] = 16'hffff;
    ctm[191] = 16'hffff;
    ctm[192] = 16'hffff;
    ctm[193] = 16'hffff;
    ctm[194] = 16'hffff;
    ctm[195] = 16'hffff;
    ctm[196] = 16'hffff;
    ctm[197] = 16'hffff;
    ctm[198] = 16'hffff;
    ctm[199] = 16'hffff;
    ctm[200] = 16'hffff;
    ctm[201] = 16'h0000;
    ctm[202] = 16'h0000;
    ctm[203] = 16'h0000;
    ctm[204] = 16'h0000;
    ctm[205] = 16'h0000;
    ctm[206] = 16'h0000;
    ctm[207] = 16'h0000;
    ctm[208] = 16'h0000;
    ctm[209] = 16'h0000;
    ctm[210] = 16'h0000;
    ctm[211] = 16'h0000;
    ctm[212] = 16'h0000;
    ctm[213] = 16'h0000;
    ctm[214] = 16'h0000;
    ctm[215] = 16'h0000;
    ctm[216] = 16'h0000;
    ctm[217] = 16'h0000;
    ctm[218] = 16'h0000;
    ctm[219] = 16'h0000;
    ctm[220] = 16'h0000;
    ctm[221] = 16'h0000;
    ctm[222] = 16'h0000;
    ctm[223] = 16'h0000;
    ctm[224] = 16'h0000;
    ctm[225] = 16'h0000;
    ctm[226] = 16'h0000;
    ctm[227] = 16'h0000;
    ctm[228] = 16'h0000;
    ctm[229] = 16'h0000;
    ctm[230] = 16'h0000;
    ctm[231] = 16'h0000;
    ctm[232] = 16'h0000;
    ctm[233] = 16'h0000;
    ctm[234] = 16'h0000;
    ctm[235] = 16'h0000;
    ctm[236] = 16'h0000;
    ctm[237] = 16'h0000;
    ctm[238] = 16'h0000;
    ctm[239] = 16'h0000;
    ctm[240] = 16'h0000;
    ctm[241] = 16'h0000;
    ctm[242] = 16'h0000;
    ctm[243] = 16'h0000;
    ctm[244] = 16'h0000;
    ctm[245] = 16'h0000;
    ctm[246] = 16'h0000;
    ctm[247] = 16'h0000;
    ctm[248] = 16'h0000;
    ctm[249] = 16'h0000;
    ctm[250] = 16'h0000;
    ctm[251] = 16'h0000;
    ctm[252] = 16'h0000;
    ctm[253] = 16'h0000;
    ctm[254] = 16'h0000;
    ctm[255] = 16'h0000;
    ctm[256] = 16'h0000;
    ctm[257] = 16'h0000;
    ctm[258] = 16'h0000;
    ctm[259] = 16'h0000;
    ctm[260] = 16'h0000;
    ctm[261] = 16'h0000;
    ctm[262] = 16'h0000;
    ctm[263] = 16'h0000;
    ctm[264] = 16'h0000;
    ctm[265] = 16'h0000;
    ctm[266] = 16'h0000;
    ctm[267] = 16'h0000;
    ctm[268] = 16'h0000;
    ctm[269] = 16'h0000;
    ctm[270] = 16'h0000;
    ctm[271] = 16'h0000;
    ctm[272] = 16'h0000;
    ctm[273] = 16'h0000;
    ctm[274] = 16'h0000;
    ctm[275] = 16'h0000;
    ctm[276] = 16'h0000;
    ctm[277] = 16'h0000;
    ctm[278] = 16'h0000;
    ctm[279] = 16'h0000;
    ctm[280] = 16'h0000;
    ctm[281] = 16'h0000;
    ctm[282] = 16'h0000;
    ctm[283] = 16'h0000;
    ctm[284] = 16'h0000;
    ctm[285] = 16'h0000;
    ctm[286] = 16'h0000;
    ctm[287] = 16'h0000;
    ctm[288] = 16'h0000;
    ctm[289] = 16'h0000;
    ctm[290] = 16'h0000;
    ctm[291] = 16'h0000;
    ctm[292] = 16'h0000;
    ctm[293] = 16'h0000;
    ctm[294] = 16'h0000;
    ctm[295] = 16'h0000;
    ctm[296] = 16'h0000;
    ctm[297] = 16'h0000;
    ctm[298] = 16'h0000;
    ctm[299] = 16'h0000;
    ctm[300] = 16'h0000;
    ctm[301] = 16'h0000;
    ctm[302] = 16'h0000;
    ctm[303] = 16'h0000;
    ctm[304] = 16'h0000;
    ctm[305] = 16'h0000;
    ctm[306] = 16'h0000;
    ctm[307] = 16'h0000;
    ctm[308] = 16'h0000;
    ctm[309] = 16'h0000;
    ctm[310] = 16'h0000;
    ctm[311] = 16'h0000;
    ctm[312] = 16'h0000;
    ctm[313] = 16'h0000;
    ctm[314] = 16'h0000;
    ctm[315] = 16'h0000;
    ctm[316] = 16'h0000;
    ctm[317] = 16'h0000;
    ctm[318] = 16'h0000;
    ctm[319] = 16'h0000;
    ctm[320] = 16'h0000;
    ctm[321] = 16'h0000;
    ctm[322] = 16'h0000;
    ctm[323] = 16'h0000;
    ctm[324] = 16'h0000;
    ctm[325] = 16'h0000;
    ctm[326] = 16'h0000;
    ctm[327] = 16'h0000;
    ctm[328] = 16'h0000;
    ctm[329] = 16'h0000;
    ctm[330] = 16'h0000;
    ctm[331] = 16'h0000;
    ctm[332] = 16'h0000;
    ctm[333] = 16'h0000;
    ctm[334] = 16'h0000;
    ctm[335] = 16'h0000;
    ctm[336] = 16'h0000;
    ctm[337] = 16'h0000;
    ctm[338] = 16'h0000;
    ctm[339] = 16'h0000;
    ctm[340] = 16'h0000;
    ctm[341] = 16'h0000;
    ctm[342] = 16'h0000;
    ctm[343] = 16'h0000;
    ctm[344] = 16'h0000;
    ctm[345] = 16'h0000;
    ctm[346] = 16'h0000;
    ctm[347] = 16'h0000;
    ctm[348] = 16'h0000;
    ctm[349] = 16'h0000;
    ctm[350] = 16'h0000;
    ctm[351] = 16'h0000;
    ctm[352] = 16'h0000;
    ctm[353] = 16'h0000;
    ctm[354] = 16'h0000;
    ctm[355] = 16'h0000;
    ctm[356] = 16'h0000;
    ctm[357] = 16'h0000;
    ctm[358] = 16'h0000;
    ctm[359] = 16'h0000;
    ctm[360] = 16'h0000;
    ctm[361] = 16'h0000;
    ctm[362] = 16'h0000;
    ctm[363] = 16'h0000;
    ctm[364] = 16'h0000;
    ctm[365] = 16'h0000;
    ctm[366] = 16'h0000;
    ctm[367] = 16'h0000;
    ctm[368] = 16'h0000;
    ctm[369] = 16'h0000;
    ctm[370] = 16'h0000;
    ctm[371] = 16'h0000;
    ctm[372] = 16'h0000;
    ctm[373] = 16'h0000;
    ctm[374] = 16'h0000;
    ctm[375] = 16'h0000;
    ctm[376] = 16'h0000;
    ctm[377] = 16'h0000;
    ctm[378] = 16'h0000;
    ctm[379] = 16'h0000;
    ctm[380] = 16'h0000;
    ctm[381] = 16'h0000;
    ctm[382] = 16'h0000;
    ctm[383] = 16'h0000;
    ctm[384] = 16'h0000;
    ctm[385] = 16'h0000;
    ctm[386] = 16'h0000;
    ctm[387] = 16'h0000;
    ctm[388] = 16'h0000;
    ctm[389] = 16'h0000;
    ctm[390] = 16'h0000;
    ctm[391] = 16'h0000;
    ctm[392] = 16'h0000;
    ctm[393] = 16'h0000;
    ctm[394] = 16'h0000;
    ctm[395] = 16'h0000;
    ctm[396] = 16'h405f;
    ctm[397] = 16'hc05f;
    ctm[398] = 16'h0000;
    ctm[399] = 16'h0000;
    ctm[400] = 16'h0000;
end
endtask

task initial_message;
begin
    message[  0] = No_Err;
    message[  1] = Res_busy;
    message[  2] = No_Food;
    message[  3] = Res_busy;
    message[  4] = No_Food;
    message[  5] = Res_busy;
    message[  6] = No_Food;
    message[  7] = Res_busy;
    message[  8] = No_Food;
    message[  9] = Res_busy;
    message[ 10] = No_Food;
    message[ 11] = Res_busy;
    message[ 12] = No_Food;
    message[ 13] = Res_busy;
    message[ 14] = No_Food;
    message[ 15] = Res_busy;
    message[ 16] = No_Food;
    message[ 17] = Res_busy;
    message[ 18] = No_Food;
    message[ 19] = Res_busy;
    message[ 20] = No_Food;
    message[ 21] = Res_busy;
    message[ 22] = Wrong_cancel;
    message[ 23] = Res_busy;
    message[ 24] = Wrong_cancel;
    message[ 25] = Res_busy;
    message[ 26] = Wrong_cancel;
    message[ 27] = Res_busy;
    message[ 28] = Wrong_cancel;
    message[ 29] = Res_busy;
    message[ 30] = Wrong_cancel;
    message[ 31] = Res_busy;
    message[ 32] = Wrong_cancel;
    message[ 33] = Res_busy;
    message[ 34] = Wrong_cancel;
    message[ 35] = Res_busy;
    message[ 36] = Wrong_cancel;
    message[ 37] = Res_busy;
    message[ 38] = Wrong_cancel;
    message[ 39] = Res_busy;
    message[ 40] = Wrong_cancel;
    message[ 41] = Res_busy;
    message[ 42] = No_customers;
    message[ 43] = Res_busy;
    message[ 44] = No_customers;
    message[ 45] = Res_busy;
    message[ 46] = No_customers;
    message[ 47] = Res_busy;
    message[ 48] = No_customers;
    message[ 49] = Res_busy;
    message[ 50] = No_customers;
    message[ 51] = Res_busy;
    message[ 52] = No_customers;
    message[ 53] = Res_busy;
    message[ 54] = No_customers;
    message[ 55] = Res_busy;
    message[ 56] = No_customers;
    message[ 57] = Res_busy;
    message[ 58] = No_customers;
    message[ 59] = Res_busy;
    message[ 60] = No_customers;
    message[ 61] = No_Food;
    message[ 62] = No_customers;
    message[ 63] = No_Food;
    message[ 64] = No_customers;
    message[ 65] = No_Food;
    message[ 66] = No_customers;
    message[ 67] = No_Food;
    message[ 68] = No_customers;
    message[ 69] = No_Food;
    message[ 70] = No_customers;
    message[ 71] = No_Food;
    message[ 72] = No_customers;
    message[ 73] = No_Food;
    message[ 74] = No_customers;
    message[ 75] = No_Food;
    message[ 76] = No_customers;
    message[ 77] = No_Food;
    message[ 78] = No_customers;
    message[ 79] = No_Food;
    message[ 80] = No_customers;
    message[ 81] = Wrong_cancel;
    message[ 82] = No_customers;
    message[ 83] = Wrong_cancel;
    message[ 84] = No_customers;
    message[ 85] = Wrong_cancel;
    message[ 86] = No_customers;
    message[ 87] = Wrong_cancel;
    message[ 88] = No_customers;
    message[ 89] = Wrong_cancel;
    message[ 90] = No_customers;
    message[ 91] = Wrong_cancel;
    message[ 92] = No_customers;
    message[ 93] = Wrong_cancel;
    message[ 94] = No_customers;
    message[ 95] = Wrong_cancel;
    message[ 96] = No_customers;
    message[ 97] = Wrong_cancel;
    message[ 98] = No_customers;
    message[ 99] = Wrong_cancel;
    message[100] = No_customers;
    message[101] = No_customers;
    message[102] = No_customers;
    message[103] = No_customers;
    message[104] = No_customers;
    message[105] = No_customers;
    message[106] = No_customers;
    message[107] = No_customers;
    message[108] = No_customers;
    message[109] = No_customers;
    message[110] = No_customers;
    message[111] = Wrong_res_ID;
    message[112] = Wrong_res_ID;
    message[113] = Wrong_res_ID;
    message[114] = Wrong_res_ID;
    message[115] = Wrong_res_ID;
    message[116] = Wrong_res_ID;
    message[117] = Wrong_res_ID;
    message[118] = Wrong_res_ID;
    message[119] = Wrong_res_ID;
    message[120] = Wrong_res_ID;
    message[121] = Wrong_res_ID;
    message[122] = Wrong_res_ID;
    message[123] = Wrong_res_ID;
    message[124] = Wrong_res_ID;
    message[125] = Wrong_res_ID;
    message[126] = Wrong_res_ID;
    message[127] = Wrong_res_ID;
    message[128] = Wrong_res_ID;
    message[129] = Wrong_res_ID;
    message[130] = Wrong_res_ID;
    message[131] = Wrong_res_ID;
    message[132] = Wrong_res_ID;
    message[133] = Wrong_res_ID;
    message[134] = Wrong_res_ID;
    message[135] = Wrong_res_ID;
    message[136] = Wrong_res_ID;
    message[137] = Wrong_res_ID;
    message[138] = Wrong_res_ID;
    message[139] = Wrong_res_ID;
    message[140] = Wrong_res_ID;
    message[141] = Wrong_food_ID;
    message[142] = Wrong_food_ID;
    message[143] = Wrong_food_ID;
    message[144] = Wrong_food_ID;
    message[145] = Wrong_food_ID;
    message[146] = Wrong_food_ID;
    message[147] = Wrong_food_ID;
    message[148] = Wrong_food_ID;
    message[149] = Wrong_food_ID;
    message[150] = Wrong_food_ID;
    message[151] = D_man_busy;
    message[152] = Wrong_food_ID;
    message[153] = D_man_busy;
    message[154] = Wrong_food_ID;
    message[155] = D_man_busy;
    message[156] = Wrong_food_ID;
    message[157] = D_man_busy;
    message[158] = Wrong_food_ID;
    message[159] = D_man_busy;
    message[160] = Wrong_food_ID;
    message[161] = D_man_busy;
    message[162] = Wrong_food_ID;
    message[163] = D_man_busy;
    message[164] = Wrong_food_ID;
    message[165] = D_man_busy;
    message[166] = Wrong_food_ID;
    message[167] = D_man_busy;
    message[168] = Wrong_food_ID;
    message[169] = D_man_busy;
    message[170] = Wrong_food_ID;
    message[171] = D_man_busy;
    message[172] = D_man_busy;
    message[173] = D_man_busy;
    message[174] = D_man_busy;
    message[175] = D_man_busy;
    message[176] = D_man_busy;
    message[177] = D_man_busy;
    message[178] = D_man_busy;
    message[179] = D_man_busy;
    message[180] = D_man_busy;
    message[181] = D_man_busy;
    message[182] = D_man_busy;
    message[183] = D_man_busy;
    message[184] = D_man_busy;
    message[185] = D_man_busy;
    message[186] = D_man_busy;
    message[187] = D_man_busy;
    message[188] = D_man_busy;
    message[189] = D_man_busy;
    message[190] = D_man_busy;
    message[191] = D_man_busy;
    message[192] = D_man_busy;
    message[193] = D_man_busy;
    message[194] = D_man_busy;
    message[195] = D_man_busy;
    message[196] = D_man_busy;
    message[197] = D_man_busy;
    message[198] = D_man_busy;
    message[199] = D_man_busy;
    message[200] = D_man_busy;
    message[201] = No_Err;
    message[202] = No_Err;
    message[203] = No_Err;
    message[204] = No_Err;
    message[205] = No_Err;
    message[206] = No_Err;
    message[207] = No_Err;
    message[208] = No_Err;
    message[209] = No_Err;
    message[210] = No_Err;
    message[211] = No_Err;
    message[212] = No_Err;
    message[213] = No_Err;
    message[214] = No_Err;
    message[215] = No_Err;
    message[216] = No_Err;
    message[217] = No_Err;
    message[218] = No_Err;
    message[219] = No_Err;
    message[220] = No_Err;
    message[221] = No_Err;
    message[222] = No_Err;
    message[223] = No_Err;
    message[224] = No_Err;
    message[225] = No_Err;
    message[226] = No_Err;
    message[227] = No_Err;
    message[228] = No_Err;
    message[229] = No_Err;
    message[230] = No_Err;
    message[231] = No_Err;
    message[232] = No_Err;
    message[233] = No_Err;
    message[234] = No_Err;
    message[235] = No_Err;
    message[236] = No_Err;
    message[237] = No_Err;
    message[238] = No_Err;
    message[239] = No_Err;
    message[240] = No_Err;
    message[241] = No_Err;
    message[242] = No_Err;
    message[243] = No_Err;
    message[244] = No_Err;
    message[245] = No_Err;
    message[246] = No_Err;
    message[247] = No_Err;
    message[248] = No_Err;
    message[249] = No_Err;
    message[250] = No_Err;
    message[251] = No_Err;
    message[252] = No_Err;
    message[253] = No_Err;
    message[254] = No_Err;
    message[255] = No_Err;
    message[256] = No_Err;
    message[257] = No_Err;
    message[258] = No_Err;
    message[259] = No_Err;
    message[260] = No_Err;
    message[261] = No_Err;
    message[262] = No_Err;
    message[263] = No_Err;
    message[264] = No_Err;
    message[265] = No_Err;
    message[266] = No_Err;
    message[267] = No_Err;
    message[268] = No_Err;
    message[269] = No_Err;
    message[270] = No_Err;
    message[271] = No_Err;
    message[272] = No_Err;
    message[273] = No_Err;
    message[274] = No_Err;
    message[275] = No_Err;
    message[276] = No_Err;
    message[277] = No_Err;
    message[278] = No_Err;
    message[279] = No_Err;
    message[280] = No_Err;
    message[281] = No_Err;
    message[282] = No_Err;
    message[283] = No_Err;
    message[284] = No_Err;
    message[285] = No_Err;
    message[286] = No_Err;
    message[287] = No_Err;
    message[288] = No_Err;
    message[289] = No_Err;
    message[290] = No_Err;
    message[291] = No_Err;
    message[292] = No_Err;
    message[293] = No_Err;
    message[294] = No_Err;
    message[295] = No_Err;
    message[296] = No_Err;
    message[297] = No_Err;
    message[298] = No_Err;
    message[299] = No_Err;
    message[300] = No_Err;
    message[301] = No_Err;
    message[302] = No_Err;
    message[303] = No_Err;
    message[304] = No_Err;
    message[305] = No_Err;
    message[306] = No_Err;
    message[307] = No_Err;
    message[308] = No_Err;
    message[309] = No_Err;
    message[310] = No_Err;
    message[311] = No_Err;
    message[312] = No_Err;
    message[313] = No_Err;
    message[314] = No_Err;
    message[315] = No_Err;
    message[316] = No_Err;
    message[317] = No_Err;
    message[318] = No_Err;
    message[319] = No_Err;
    message[320] = No_Err;
    message[321] = No_Err;
    message[322] = No_Err;
    message[323] = No_Err;
    message[324] = No_Err;
    message[325] = No_Err;
    message[326] = No_Err;
    message[327] = No_Err;
    message[328] = No_Err;
    message[329] = No_Err;
    message[330] = No_Err;
    message[331] = No_Err;
    message[332] = No_Err;
    message[333] = No_Err;
    message[334] = No_Err;
    message[335] = No_Err;
    message[336] = No_Err;
    message[337] = No_Err;
    message[338] = No_Err;
    message[339] = No_Err;
    message[340] = No_Err;
    message[341] = No_Err;
    message[342] = No_Err;
    message[343] = No_Err;
    message[344] = No_Err;
    message[345] = No_Err;
    message[346] = No_Err;
    message[347] = No_Err;
    message[348] = No_Err;
    message[349] = No_Err;
    message[350] = No_Err;
    message[351] = No_Err;
    message[352] = No_Err;
    message[353] = No_Err;
    message[354] = No_Err;
    message[355] = No_Err;
    message[356] = No_Err;
    message[357] = No_Err;
    message[358] = No_Err;
    message[359] = No_Err;
    message[360] = No_Err;
    message[361] = No_Err;
    message[362] = No_Err;
    message[363] = No_Err;
    message[364] = No_Err;
    message[365] = No_Err;
    message[366] = No_Err;
    message[367] = No_Err;
    message[368] = No_Err;
    message[369] = No_Err;
    message[370] = No_Err;
    message[371] = No_Err;
    message[372] = No_Err;
    message[373] = No_Err;
    message[374] = No_Err;
    message[375] = No_Err;
    message[376] = No_Err;
    message[377] = No_Err;
    message[378] = No_Err;
    message[379] = No_Err;
    message[380] = No_Err;
    message[381] = No_Err;
    message[382] = No_Err;
    message[383] = No_Err;
    message[384] = No_Err;
    message[385] = No_Err;
    message[386] = No_Err;
    message[387] = No_Err;
    message[388] = No_Err;
    message[389] = No_Err;
    message[390] = No_Err;
    message[391] = No_Err;
    message[392] = No_Err;
    message[393] = No_Err;
    message[394] = No_Err;
    message[395] = No_Err;
    message[396] = No_Err;
    message[397] = No_Err;
    message[398] = No_Err;
    message[399] = No_Err;
    message[400] = No_Err;
end
endtask

task initial_answer;
begin
    answer[  0] = 64'b0;
    answer[  1] = 64'b0;
    answer[  2] = 64'b0;
    answer[  3] = 64'b0;
    answer[  4] = 64'b0;
    answer[  5] = 64'b0;
    answer[  6] = 64'b0;
    answer[  7] = 64'b0;
    answer[  8] = 64'b0;
    answer[  9] = 64'b0;
    answer[ 10] = 64'b0;
    answer[ 11] = 64'b0;
    answer[ 12] = 64'b0;
    answer[ 13] = 64'b0;
    answer[ 14] = 64'b0;
    answer[ 15] = 64'b0;
    answer[ 16] = 64'b0;
    answer[ 17] = 64'b0;
    answer[ 18] = 64'b0;
    answer[ 19] = 64'b0;
    answer[ 20] = 64'b0;
    answer[ 21] = 64'b0;
    answer[ 22] = 64'b0;
    answer[ 23] = 64'b0;
    answer[ 24] = 64'b0;
    answer[ 25] = 64'b0;
    answer[ 26] = 64'b0;
    answer[ 27] = 64'b0;
    answer[ 28] = 64'b0;
    answer[ 29] = 64'b0;
    answer[ 30] = 64'b0;
    answer[ 31] = 64'b0;
    answer[ 32] = 64'b0;
    answer[ 33] = 64'b0;
    answer[ 34] = 64'b0;
    answer[ 35] = 64'b0;
    answer[ 36] = 64'b0;
    answer[ 37] = 64'b0;
    answer[ 38] = 64'b0;
    answer[ 39] = 64'b0;
    answer[ 40] = 64'b0;
    answer[ 41] = 64'b0;
    answer[ 42] = 64'b0;
    answer[ 43] = 64'b0;
    answer[ 44] = 64'b0;
    answer[ 45] = 64'b0;
    answer[ 46] = 64'b0;
    answer[ 47] = 64'b0;
    answer[ 48] = 64'b0;
    answer[ 49] = 64'b0;
    answer[ 50] = 64'b0;
    answer[ 51] = 64'b0;
    answer[ 52] = 64'b0;
    answer[ 53] = 64'b0;
    answer[ 54] = 64'b0;
    answer[ 55] = 64'b0;
    answer[ 56] = 64'b0;
    answer[ 57] = 64'b0;
    answer[ 58] = 64'b0;
    answer[ 59] = 64'b0;
    answer[ 60] = 64'b0;
    answer[ 61] = 64'b0;
    answer[ 62] = 64'b0;
    answer[ 63] = 64'b0;
    answer[ 64] = 64'b0;
    answer[ 65] = 64'b0;
    answer[ 66] = 64'b0;
    answer[ 67] = 64'b0;
    answer[ 68] = 64'b0;
    answer[ 69] = 64'b0;
    answer[ 70] = 64'b0;
    answer[ 71] = 64'b0;
    answer[ 72] = 64'b0;
    answer[ 73] = 64'b0;
    answer[ 74] = 64'b0;
    answer[ 75] = 64'b0;
    answer[ 76] = 64'b0;
    answer[ 77] = 64'b0;
    answer[ 78] = 64'b0;
    answer[ 79] = 64'b0;
    answer[ 80] = 64'b0;
    answer[ 81] = 64'b0;
    answer[ 82] = 64'b0;
    answer[ 83] = 64'b0;
    answer[ 84] = 64'b0;
    answer[ 85] = 64'b0;
    answer[ 86] = 64'b0;
    answer[ 87] = 64'b0;
    answer[ 88] = 64'b0;
    answer[ 89] = 64'b0;
    answer[ 90] = 64'b0;
    answer[ 91] = 64'b0;
    answer[ 92] = 64'b0;
    answer[ 93] = 64'b0;
    answer[ 94] = 64'b0;
    answer[ 95] = 64'b0;
    answer[ 96] = 64'b0;
    answer[ 97] = 64'b0;
    answer[ 98] = 64'b0;
    answer[ 99] = 64'b0;
    answer[100] = 64'b0;
    answer[101] = 64'b0;
    answer[102] = 64'b0;
    answer[103] = 64'b0;
    answer[104] = 64'b0;
    answer[105] = 64'b0;
    answer[106] = 64'b0;
    answer[107] = 64'b0;
    answer[108] = 64'b0;
    answer[109] = 64'b0;
    answer[110] = 64'b0;
    answer[111] = 64'b0;
    answer[112] = 64'b0;
    answer[113] = 64'b0;
    answer[114] = 64'b0;
    answer[115] = 64'b0;
    answer[116] = 64'b0;
    answer[117] = 64'b0;
    answer[118] = 64'b0;
    answer[119] = 64'b0;
    answer[120] = 64'b0;
    answer[121] = 64'b0;
    answer[122] = 64'b0;
    answer[123] = 64'b0;
    answer[124] = 64'b0;
    answer[125] = 64'b0;
    answer[126] = 64'b0;
    answer[127] = 64'b0;
    answer[128] = 64'b0;
    answer[129] = 64'b0;
    answer[130] = 64'b0;
    answer[131] = 64'b0;
    answer[132] = 64'b0;
    answer[133] = 64'b0;
    answer[134] = 64'b0;
    answer[135] = 64'b0;
    answer[136] = 64'b0;
    answer[137] = 64'b0;
    answer[138] = 64'b0;
    answer[139] = 64'b0;
    answer[140] = 64'b0;
    answer[141] = 64'b0;
    answer[142] = 64'b0;
    answer[143] = 64'b0;
    answer[144] = 64'b0;
    answer[145] = 64'b0;
    answer[146] = 64'b0;
    answer[147] = 64'b0;
    answer[148] = 64'b0;
    answer[149] = 64'b0;
    answer[150] = 64'b0;
    answer[151] = 64'b0;
    answer[152] = 64'b0;
    answer[153] = 64'b0;
    answer[154] = 64'b0;
    answer[155] = 64'b0;
    answer[156] = 64'b0;
    answer[157] = 64'b0;
    answer[158] = 64'b0;
    answer[159] = 64'b0;
    answer[160] = 64'b0;
    answer[161] = 64'b0;
    answer[162] = 64'b0;
    answer[163] = 64'b0;
    answer[164] = 64'b0;
    answer[165] = 64'b0;
    answer[166] = 64'b0;
    answer[167] = 64'b0;
    answer[168] = 64'b0;
    answer[169] = 64'b0;
    answer[170] = 64'b0;
    answer[171] = 64'b0;
    answer[172] = 64'b0;
    answer[173] = 64'b0;
    answer[174] = 64'b0;
    answer[175] = 64'b0;
    answer[176] = 64'b0;
    answer[177] = 64'b0;
    answer[178] = 64'b0;
    answer[179] = 64'b0;
    answer[180] = 64'b0;
    answer[181] = 64'b0;
    answer[182] = 64'b0;
    answer[183] = 64'b0;
    answer[184] = 64'b0;
    answer[185] = 64'b0;
    answer[186] = 64'b0;
    answer[187] = 64'b0;
    answer[188] = 64'b0;
    answer[189] = 64'b0;
    answer[190] = 64'b0;
    answer[191] = 64'b0;
    answer[192] = 64'b0;
    answer[193] = 64'b0;
    answer[194] = 64'b0;
    answer[195] = 64'b0;
    answer[196] = 64'b0;
    answer[197] = 64'b0;
    answer[198] = 64'b0;
    answer[199] = 64'b0;
    answer[200] = 64'b0;
    answer[201] = {16'hffff, 48'b0};
    answer[202] = 64'b0;
    answer[203] = 64'b0;
    answer[204] = 64'b0;
    answer[205] = 64'b0;
    answer[206] = 64'b0;
    answer[207] = 64'b0;
    answer[208] = 64'b0;
    answer[209] = 64'b0;
    answer[210] = 64'b0;
    answer[211] = 64'b0;
    answer[212] = 64'b0;
    answer[213] = 64'b0;
    answer[214] = 64'b0;
    answer[215] = 64'b0;
    answer[216] = 64'b0;
    answer[217] = 64'b0;
    answer[218] = 64'b0;
    answer[219] = 64'b0;
    answer[220] = 64'b0;
    answer[221] = 64'b0;
    answer[222] = 64'b0;
    answer[223] = 64'b0;
    answer[224] = 64'b0;
    answer[225] = 64'b0;
    answer[226] = 64'b0;
    answer[227] = 64'b0;
    answer[228] = 64'b0;
    answer[229] = 64'b0;
    answer[230] = 64'b0;
    answer[231] = 64'b0;
    answer[232] = 64'b0;
    answer[233] = 64'b0;
    answer[234] = 64'b0;
    answer[235] = 64'b0;
    answer[236] = 64'b0;
    answer[237] = 64'b0;
    answer[238] = 64'b0;
    answer[239] = 64'b0;
    answer[240] = 64'b0;
    answer[241] = 64'b0;
    answer[242] = 64'b0;
    answer[243] = 64'b0;
    answer[244] = 64'b0;
    answer[245] = 64'b0;
    answer[246] = 64'b0;
    answer[247] = 64'b0;
    answer[248] = 64'b0;
    answer[249] = 64'b0;
    answer[250] = 64'b0;
    answer[251] = 64'b0;
    answer[252] = 64'b0;
    answer[253] = 64'b0;
    answer[254] = 64'b0;
    answer[255] = 64'b0;
    answer[256] = 64'b0;
    answer[257] = 64'b0;
    answer[258] = 64'b0;
    answer[259] = 64'b0;
    answer[260] = 64'b0;
    answer[261] = 64'b0;
    answer[262] = 64'b0;
    answer[263] = 64'b0;
    answer[264] = 64'b0;
    answer[265] = 64'b0;
    answer[266] = 64'b0;
    answer[267] = 64'b0;
    answer[268] = 64'b0;
    answer[269] = 64'b0;
    answer[270] = 64'b0;
    answer[271] = 64'b0;
    answer[272] = 64'b0;
    answer[273] = 64'b0;
    answer[274] = 64'b0;
    answer[275] = 64'b0;
    answer[276] = 64'b0;
    answer[277] = 64'b0;
    answer[278] = 64'b0;
    answer[279] = 64'b0;
    answer[280] = 64'b0;
    answer[281] = 64'b0;
    answer[282] = 64'b0;
    answer[283] = 64'b0;
    answer[284] = 64'b0;
    answer[285] = 64'b0;
    answer[286] = 64'b0;
    answer[287] = 64'hfd030100;
    answer[288] = 64'hfd040100;
    answer[289] = 64'hfd050100;
    answer[290] = 64'hfd060100;
    answer[291] = 64'hfd070100;
    answer[292] = 64'hfd080100;
    answer[293] = 64'hfd090100;
    answer[294] = 64'hfd0a0100;
    answer[295] = 64'hfd0b0100;
    answer[296] = 64'hfd0c0100;
    answer[297] = 64'hfd0d0100;
    answer[298] = 64'hfd0e0100;
    answer[299] = 64'hfd0f0100;
    answer[300] = 64'hfd100100;
    answer[301] = 64'hfd110100;
    answer[302] = 64'hfd120100;
    answer[303] = 64'hfd130100;
    answer[304] = 64'hfd140100;
    answer[305] = 64'hfd150100;
    answer[306] = 64'hfd160100;
    answer[307] = 64'hfd170100;
    answer[308] = 64'hfd180100;
    answer[309] = 64'hfd190100;
    answer[310] = 64'hfd1a0100;
    answer[311] = 64'hfd1b0100;
    answer[312] = 64'hfd1c0100;
    answer[313] = 64'hfd1d0100;
    answer[314] = 64'hfd1e0100;
    answer[315] = 64'hfd1f0100;
    answer[316] = 64'hfd200100;
    answer[317] = 64'hfd210100;
    answer[318] = 64'hfd220100;
    answer[319] = 64'hfd230100;
    answer[320] = 64'hfd240100;
    answer[321] = 64'hfd250100;
    answer[322] = 64'hfd260100;
    answer[323] = 64'hfd270100;
    answer[324] = 64'hfd280100;
    answer[325] = 64'hfd290100;
    answer[326] = 64'hfd2a0100;
    answer[327] = 64'hfd2b0100;
    answer[328] = 64'hfd2c0100;
    answer[329] = 64'hfd2d0100;
    answer[330] = 64'hfd2e0100;
    answer[331] = 64'hfd2f0100;
    answer[332] = 64'hfd300100;
    answer[333] = 64'hfd310100;
    answer[334] = 64'hfd320100;
    answer[335] = 64'hfd330100;
    answer[336] = 64'hfd340100;
    answer[337] = 64'hfd350100;
    answer[338] = 64'hfd360100;
    answer[339] = 64'hfd370100;
    answer[340] = 64'hfd380100;
    answer[341] = 64'hfd390100;
    answer[342] = 64'hfd3a0100;
    answer[343] = 64'hfd3b0100;
    answer[344] = 64'hfd3c0100;
    answer[345] = 64'hfd3d0100;
    answer[346] = 64'hfd3e0100;
    answer[347] = 64'hfd3f0100;
    answer[348] = 64'hfd400100;
    answer[349] = 64'hfd410100;
    answer[350] = 64'hfd420100;
    answer[351] = 64'hfd430100;
    answer[352] = 64'hfd440100;
    answer[353] = 64'hfd450100;
    answer[354] = 64'hfd460100;
    answer[355] = 64'hfd470100;
    answer[356] = 64'hfd480100;
    answer[357] = 64'hfd490100;
    answer[358] = 64'hfd4a0100;
    answer[359] = 64'hfd4b0100;
    answer[360] = 64'hfd4c0100;
    answer[361] = 64'hfd4d0100;
    answer[362] = 64'hfd4e0100;
    answer[363] = 64'hfd4f0100;
    answer[364] = 64'hfd500100;
    answer[365] = 64'hfd510100;
    answer[366] = 64'hfd520100;
    answer[367] = 64'hfd530100;
    answer[368] = 64'hfd540100;
    answer[369] = 64'hfd550100;
    answer[370] = 64'hfd560100;
    answer[371] = 64'hfd570100;
    answer[372] = 64'hfd580100;
    answer[373] = 64'hfd590100;
    answer[374] = 64'hfd5a0100;
    answer[375] = 64'hfd5b0100;
    answer[376] = 64'hfd5c0100;
    answer[377] = 64'hfd5d0100;
    answer[378] = 64'hfd5e0100;
    answer[379] = 64'hfd5f0100;
    answer[380] = 64'hfd600100;
    answer[381] = 64'hfd610100;
    answer[382] = 64'hfd620100;
    answer[383] = 64'hfd630100;
    answer[384] = 64'hfd640100;
    answer[385] = 64'hfd650100;
    answer[386] = 64'hfd660100;
    answer[387] = 64'hfd670100;
    answer[388] = 64'hfd680100;
    answer[389] = 64'hfd690100;
    answer[390] = 64'hfd6a0100;
    answer[391] = 64'hfd6b0100;
    answer[392] = 64'hfd6c0100;
    answer[393] = 64'hfd6d0100;
    answer[394] = 64'hfd6e0100;
    answer[395] = {16'hfdff, 48'b0};
    answer[396] = {16'h405f, 16'b0, 32'hfd404f4f};
    answer[397] = {32'hc05f405f, 32'hfd314f4f};
    answer[398] = 64'b0;
    answer[399] = {16'hfdff, 48'b0};
    answer[400] = 64'b0;
end
endtask

endprogram
